//////////////////////////////////////
///T.Guru Nandini Devi             ///
///nandinidevitekumudi@gmail.com   ///
///Submission Date: 25-07-2025     ///
//////////////////////////////////////
//Implement the wire circuit
module top_module (
    input in,
    output out);
   assign out = in;
endmodule


