//////////////////////////////////////
///T.Guru Nandini Devi             ///
///nandinidevitekumudi@gmail.com   ///
///Submission Date: 26-05-2025     ///
//////////////////////////////////////
//Create a module that implements an AND gate.
module top_module( 
    input a, 
    input b, 
    output out );
    assign out = a & b;
endmodule
