////////////////////////////////////////
// T.Guru Nandini Devi
// nandinidevitekumudi@gmail.com
// submission date: 21-05-2025
/////////////////////////////////////////
//Problem Statement - 02 : Build a circuit with no inputs and one output that outputs a constant 0
module top_module(
    output zero
);
  // Module body starts after semicolon
assign zero=1'b0;
endmodule
