//////////////////////////////////////
///T.Guru Nandini Devi             ///
///nandinidevitekumudi@gmail.com   ///
///Submission Date: 22-05-2025     ///
//////////////////////////////////////
//Create a module that implements a NOT gate.
module top_module(
  input in, 
  output out 
);
assign out= ~in;
endmodule
