//////////////////////////////////////
///T.Guru Nandini Devi             ///
///nandinidevitekumudi@gmail.com   ///
//////////////////////////////////////
//Implement Ground circuit
module top_module (
    output out);
   assign out=1'b0;
endmodule
