////////////////////////////////////////
// T.Guru Nandini Devi
// nandinidevitekumudi@gmail.com
// submission date: 20-05-2025
/////////////////////////////////////////
//Build a circuit with no inputs and one output. That output should always drive 1 (or logic high).
module top_module( output one );

// Insert your code here
    assign one = 1'b1;

endmodule
